module image

//
