module viup

struct Control {
	ptr      voidptr
	@type    string
}