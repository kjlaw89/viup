module viup

pub enum Pos {
	center       = 0xFFFF
	left         = 0xFFFE
	right        = 0xFFFD
	mousepos     = 0xFFFC
	current      = 0xFFFB
	centerparent = 0xFFFA
	leftparent   = 0xFFF9
	rightparent  = 0xFFF8
}