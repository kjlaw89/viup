module image

// 